//ALU
`include "PCPU_ctrl_encode_def.v"

module alu(A, B, ALUOp, C, Zero);
           
   input  signed [31:0] A, B;
   input         [3:0]  ALUOp;
   output signed [31:0] C;
   output Zero;
   
   reg [31:0] C_temp;
   reg [31:0] C;
   
   always @( A or B or ALUOp ) begin    ///////////////////////////////////changed
      case ( ALUOp )
          `ALU_NOP:  C = A;                          // NOP
          `ALU_ADD:  C = A + B;                      // ADD/ADDI
          `ALU_ADDU: C = A + B;                      // ADDU
          `ALU_SUBU: C = A - B;                      // SUBU
          `ALU_SUB:  C = A - B;                      // SUB
          `ALU_AND:  C = A & B;                      // AND/ANDI
          `ALU_OR:   C = A | B;                      // OR/ORI
          `ALU_SLT:  C = (A < B) ? 32'd1 : 32'd0;    // SLT/SLTI
          `ALU_SLTU: C = ({1'b0, A} < {1'b0, B}) ? 32'd1 : 32'd0;//SLTU
          `ALU_NOR:  C = ~(A | B);                   //NOR
          `ALU_LUI:  C = {B[15:0],16'b0};            //LUI
          default:   C = A;                          // Undefined
      endcase
   end // end always
   
   assign Zero = (C == 32'b0);

endmodule
    
